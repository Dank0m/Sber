module  blackbox            // module - ключевое слово, blackbox - имя модуля
#(
                            //Здесь могут находиться параметры
)
(
    input  a, b, c          // входные порты a,b,c
    input  [7:0] bus,       // входной порт bus - 8-разрядная шина
    output  [7:0] bus_out   // выходной порт bus_out, также 8-разрядный
);
                            // Здесь добавляется тело модуля

endmodule                   // endmodule - конец описания модуля, ключевое слово
