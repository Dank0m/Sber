`timescale 1ns / 100ps

module testbench();
    // Тактовый генератор
    reg clk = 1'b0;
    always begin
        #5 clk = ~clk;  // Инверсия каждые 5 наносекунд
    end
    // Входной сигнал для подключения к тестируемому модулю
    reg signal_i = 1'b0;
    // Выходной сигнал для подключения к тестируемому модулю
    wire signal_o;
    
    // Экземпляр тестируемого модуля
    overlay imported_module(
//синтаксис: module_name instance_name
/*module_name — Имя модуля которое даем модулю при его объявлении*/
/*instance_name — Имя экземпляра. Это уникальное имя, которое вы 
даете конкретному экземпляру модуля, когда используете его в 
другом модуле или тестбенче.*/
        .clk_i(clk), 
        .a_i(signal_i),
        .a_o(signal_o)
//синтаксис: .порт_модуля_который_тестируем(порт_который_описан_в_testbench)
    );
    
    // Блок инициализации
    initial begin
        $dumpvars;
        #10; 
        signal_i <= ~signal_i;
        #10; 
        signal_i <= ~signal_i;
        #10; 
        signal_i <= ~signal_i;
        #10;                          
        $finish;                      // Завершение симуляции
    end
    /*Initial — это процедурный блок, который описывает поведение 
    в начале симуляции. Он позволяет инициализировать переменные и
    задавать конкретные значения портам дизайна в начале моделирования.
    Выполнение начального блока начинается в момент времени 0 в 
    симуляции. Он выполняется только один раз во время симуляции и 
    завершается, когда выполнены все содержащиеся в нём операторы
    */
endmodule
